
`define rows        6
`define cols        4
`define AW          20
`define DW          32
`define CFGW        (`AW + `DW)
`define CFG_LENGTH  133